* On-die Decoupling circuit for z11b (VDDQ to VSSQ)
* Includes VDDQ-VSSQ decoupling for an individual signal such as DQ0-15, LDQS_t/c, UDQS_t/c, UDM or LDM.
* This subcircuit should be added across the IBIS DQ, DM or DQS model's [Pullup Reference] and [Pulldown Reference]
* nodes as in the following Spice example:

******************************************************************************************************
*x_decouple vddq_die vss_die gnd z11b_ondie_decoupling_perdq

*b_dq1 vccq_die vss_die PAD_DQ1 IN_DQ1 ENOUT RCVR_OUT_DQ1 vccq_die vss_die
*+ file='z11b.ibs' model='DQ_34_2933' typ=typ power=off buffer=3 interpol=1 ramp_fwf=2 ramp_rwf=2
*+ rm_tail_rwf=default rm_tail_fwf=default
*+ rm_dly_rwf=default rm_dly_fwf=default
******************************************************************************************************

.subckt z11b_ondie_decoupling_perdq vddq_die vss_die ref
x1 vddq_die vss_die ref cfat_perdq_sparam_50

**********************************************************
** STATE-SPACE REALIZATION
** IN SPICE LANGUAGE
** This file is automatically generated
**********************************************************
** Created: 23-Aug-2019 by IdEM MP 12 (12.1.0)
**********************************************************
**
**********************************************************
** COMMENTS
**********************************************************
**
**  NPort=2 DATA=1332 NOISE=0 GROUPDELAY=0 COMPLEX_DATAFORMAT=POLAR
**  NumOfBlock=1 NumOfParam=0
** 
**  .MODEL Smodel S TSTONEFILE=cfat_perdq_sparam_50.s2p TYPE=S
**    -- The above .MODEL line can be used for the S element in the netlist.
** 
** 
**
**********************************************************
**
**
**---------------------------
** Options Used in IdEM Flow
**---------------------------
**
** Fitting Options **
**
** Bandwidth: 2.0417e+10 Hz
** Order: [2 2 6] 
** SplitType: none 
** tol: 1.0000e-04 
**
**---------------------------
**
** Passivity Options **
**
** Alg: SOC+HAM 
**    Max SOC it: 50 
**    Max HAM it: 50 
** Freq sampling: manual
**    In-band samples: 200
**    Off-band samples: 100
** Optimization method: Model based
**
**---------------------------
**
** Netlist Options **
**
** Netlist format: SPICE standard
** Port reference: common
** Voltage-controlled current sources
**
**---------------------------
**
**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* ref  --> reference node, common for all the input nodes 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt cfat_perdq_sparam_50
+  a_1 a_2 ref
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
GRI_1 NI_1 ref NI_1 ref 2.0000000000000000e-02
GC_1_1 ref NI_1 NS_1 0 7.5822795216346096e-03
GC_1_2 ref NI_1 NS_2 0 3.5902013174278755e-03
GC_1_3 ref NI_1 NS_3 0 7.2846812529359624e-03
GC_1_4 ref NI_1 NS_4 0 3.1695903643706329e-02
GC_1_5 ref NI_1 NS_5 0 5.4660964083090450e-07
GC_1_6 ref NI_1 NS_6 0 1.4926463349190639e-04
GC_1_7 ref NI_1 NS_7 0 -3.6739983615024862e-04
GC_1_8 ref NI_1 NS_8 0 -4.0509249447121401e-03
GC_1_9 ref NI_1 NS_9 0 -7.2051350599292349e-03
GC_1_10 ref NI_1 NS_10 0 -3.1739261413559886e-02
GC_1_11 ref NI_1 NS_11 0 -1.1639787203465530e-06
GC_1_12 ref NI_1 NS_12 0 -1.4443429342608907e-04
GD_1_1 ref NI_1 NA_1 0 9.3536045431372398e-03
GD_1_2 ref NI_1 NA_2 0 2.7320626521876606e-01
*
* Port 2
VI_2 a_2 NI_2 0
GRI_2 NI_2 ref NI_2 ref 2.0000000000000000e-02
GC_2_1 ref NI_2 NS_1 0 -3.6739985184936456e-04
GC_2_2 ref NI_2 NS_2 0 -4.0509249438178954e-03
GC_2_3 ref NI_2 NS_3 0 -7.2051350598360498e-03
GC_2_4 ref NI_2 NS_4 0 -3.1739261413545446e-02
GC_2_5 ref NI_2 NS_5 0 -1.1639787204915532e-06
GC_2_6 ref NI_2 NS_6 0 -1.4443429341980951e-04
GC_2_7 ref NI_2 NS_7 0 7.5822795189273021e-03
GC_2_8 ref NI_2 NS_8 0 3.5902013166808403e-03
GC_2_9 ref NI_2 NS_9 0 7.2846812539232733e-03
GC_2_10 ref NI_2 NS_10 0 3.1695903643698793e-02
GC_2_11 ref NI_2 NS_11 0 5.4660963371374044e-07
GC_2_12 ref NI_2 NS_12 0 1.4926463354163091e-04
GD_2_1 ref NI_2 NA_1 0 2.7320626521857244e-01
GD_2_2 ref NI_2 NA_2 0 9.3536045438131956e-03
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
GRA_1 NA_1 0 NA_1 0 2.8284271247461901e-01
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 ref 2.0000000000000000e-02
*
* Impinging wave, port 2
GRA_2 NA_2 0 NA_2 0 2.8284271247461901e-01
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 ref 2.0000000000000000e-02
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 1.0000000000000001e-09
GRS_1 NS_1 0 NS_1 0 5.2707388993577524e+00
GS_1_1 0 NS_1 NA_1 0 2.2427717688837773e-01
*
* Real pole n. 2
CS_2 NS_2 0 1.0000000000000001e-09
GRS_2 NS_2 0 NS_2 0 7.3434129992739949e-01
GS_2_1 0 NS_2 NA_1 0 2.2427717688837773e-01
*
* Real pole n. 3
CS_3 NS_3 0 1.0000000000000001e-09
GRS_3 NS_3 0 NS_3 0 7.0517678890748836e-02
GS_3_1 0 NS_3 NA_1 0 2.2427717688837773e-01
*
* Real pole n. 4
CS_4 NS_4 0 1.0000000000000001e-09
GRS_4 NS_4 0 NS_4 0 2.9249610747441535e-02
GS_4_1 0 NS_4 NA_1 0 2.2427717688837773e-01
*
* Real pole n. 5
CS_5 NS_5 0 1.0000000000000001e-09
GRS_5 NS_5 0 NS_5 0 5.1192535935390762e-04
GS_5_1 0 NS_5 NA_1 0 2.2427717688837773e-01
*
* Real pole n. 6
CS_6 NS_6 0 1.0000000000000001e-09
GRS_6 NS_6 0 NS_6 0 6.1092836856464971e-03
GS_6_1 0 NS_6 NA_1 0 2.2427717688837773e-01
*
* Real pole n. 7
CS_7 NS_7 0 1.0000000000000001e-09
GRS_7 NS_7 0 NS_7 0 5.2707388993577524e+00
GS_7_2 0 NS_7 NA_2 0 2.2427717688837773e-01
*
* Real pole n. 8
CS_8 NS_8 0 1.0000000000000001e-09
GRS_8 NS_8 0 NS_8 0 7.3434129992739949e-01
GS_8_2 0 NS_8 NA_2 0 2.2427717688837773e-01
*
* Real pole n. 9
CS_9 NS_9 0 1.0000000000000001e-09
GRS_9 NS_9 0 NS_9 0 7.0517678890748836e-02
GS_9_2 0 NS_9 NA_2 0 2.2427717688837773e-01
*
* Real pole n. 10
CS_10 NS_10 0 1.0000000000000001e-09
GRS_10 NS_10 0 NS_10 0 2.9249610747441535e-02
GS_10_2 0 NS_10 NA_2 0 2.2427717688837773e-01
*
* Real pole n. 11
CS_11 NS_11 0 1.0000000000000001e-09
GRS_11 NS_11 0 NS_11 0 5.1192535935390762e-04
GS_11_2 0 NS_11 NA_2 0 2.2427717688837773e-01
*
* Real pole n. 12
CS_12 NS_12 0 1.0000000000000001e-09
GRS_12 NS_12 0 NS_12 0 6.1092836856464971e-03
GS_12_2 0 NS_12 NA_2 0 2.2427717688837773e-01
*
******************************


.ends
.ends
*******************
* End of subcircuit
*******************
